LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE IEEE.std_logic_unsigned.ALL;

ENTITY BRANCH_CONTROL IS
    PORT (
        CLK, RESET, HAS_NEXT_OPERAND, BRANCH, JMP : IN STD_LOGIC;
        PC_IN, R_DEST_ADDRESS : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
        OPCODE : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
        FLAGS : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
        IS_BRANCH_TAKEN : OUT STD_LOGIC;
        PC_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
END BRANCH_CONTROL;

ARCHITECTURE ARCH_BRANCH_CONTROL OF BRANCH_CONTROL IS

    SIGNAL COMPARATOR_OUT : STD_LOGIC;
    SIGNAL BRANCH_TAKEN_SIG : STD_LOGIC;
    SIGNAL ADDER_OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL FLAGS_OPCODE_CHECKER : STD_LOGIC_VECTOR(4 DOWNTO 0);

BEGIN

    PROCESS (CLK, RESET)
    BEGIN

        IF RESET = '1' THEN

            IS_BRANCH_TAKEN <= '0';
            PC_OUT <= (OTHERS => '0');

        ELSIF RISING_EDGE(CLK) THEN
            -- COMBINING THE LAST TWO BITS IN OPCODE WITH THE FLAGS BITS
            FLAGS_OPCODE_CHECKER <= OPCODE(1 DOWNTO 0) & FLAGS(2 DOWNTO 0);
            CASE FLAGS_OPCODE_CHECKER IS
                WHEN "01001" => COMPARATOR_OUT <= '1';
                WHEN "10010" => COMPARATOR_OUT <= '1';
                WHEN "11100" => COMPARATOR_OUT <= '1';
                WHEN OTHERS => COMPARATOR_OUT <= '0';
            END CASE;

            IS_BRANCH_TAKEN <= (COMPARATOR_OUT AND BRANCH) OR JMP;
            BRANCH_TAKEN_SIG <= (COMPARATOR_OUT AND BRANCH) OR JMP;

            IF HAS_NEXT_OPERAND = '1' THEN
                ADDER_OUT <= PC_IN + 4;
            ELSE
                ADDER_OUT <= PC_IN + 2;
            END IF;

            IF BRANCH_TAKEN_SIG = '1' THEN
                PC_OUT <= R_DEST_ADDRESS;
            ELSE
                PC_OUT <= ADDER_OUT;
            END IF;

        END IF;
    END PROCESS;

END ARCHITECTURE;