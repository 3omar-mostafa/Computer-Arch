LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE IEEE.std_logic_unsigned.ALL;

ENTITY BRANCH_CONTROL IS
    PORT (
        CLK, RESET, HAS_NEXT_OPERAND, BRANCH, JMP : IN STD_LOGIC;
        PC_IN, R_DEST_ADDRESS : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
        OPCODE : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
        carry_flag    : IN STD_LOGIC;
		negative_flag : IN STD_LOGIC;
		zero_flag     : IN STD_LOGIC;
        IS_BRANCH_TAKEN : OUT STD_LOGIC;
        PC_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
END BRANCH_CONTROL;

ARCHITECTURE ARCH_BRANCH_CONTROL OF BRANCH_CONTROL IS

    SIGNAL COMPARATOR_OUT : STD_LOGIC;
    SIGNAL BRANCH_TAKEN_SIG : STD_LOGIC;
    SIGNAL ADDER_OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL FLAGS_OPCODE_CHECKER : STD_LOGIC_VECTOR(4 DOWNTO 0);

BEGIN

    -- COMBINING THE LAST TWO BITS IN OPCODE WITH THE FLAGS BITS
    FLAGS_OPCODE_CHECKER <= OPCODE(1 DOWNTO 0) & carry_flag & negative_flag & zero_flag;

    COMPARATOR_OUT <= '1' WHEN (FLAGS_OPCODE_CHECKER = "01001" OR FLAGS_OPCODE_CHECKER = "10010" OR FLAGS_OPCODE_CHECKER = "11100")
                 ELSE '0';

    BRANCH_TAKEN_SIG <= (COMPARATOR_OUT AND BRANCH) OR JMP;

    ADDER_OUT <= (PC_IN + 2) WHEN HAS_NEXT_OPERAND = '1'
        ELSE (PC_IN + 1);

    PC_OUT <= R_DEST_ADDRESS WHEN BRANCH_TAKEN_SIG = '1'
         ELSE ADDER_OUT;

    PROCESS(CLK)
    BEGIN
        IF FALLING_EDGE(CLK) THEN
            IS_BRANCH_TAKEN <= '0';
        ELSIF RISING_EDGE(CLK) THEN
            IS_BRANCH_TAKEN <= BRANCH_TAKEN_SIG;
        END IF;
    END PROCESS;

END ARCHITECTURE;