LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY CONTROL_UNIT IS
	PORT (
		CLK, RESET : IN STD_LOGIC;
		IR : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		IS_LOAD_STORE, MEM_READ, MEM_WRITE, WRITE_BACK, BRANCH, JMP, HAS_NEXT_OPERAND, PUSH, POP : OUT STD_LOGIC
	);
END CONTROL_UNIT;

ARCHITECTURE ARCH_CONTROL_UNIT OF CONTROL_UNIT IS

BEGIN

	PROCESS (CLK, RESET)

	BEGIN

		IF RESET = '1' THEN

			IS_LOAD_STORE <= '0';
			MEM_READ <= '0';
			MEM_WRITE <= '0';
			WRITE_BACK <= '0';
			BRANCH <= '0';
			JMP <= '0';
			HAS_NEXT_OPERAND <= '0';
			PUSH <= '0';
			POP <= '0';

		ELSIF RISING_EDGE(CLK) THEN

			IS_LOAD_STORE <= (IR(31) AND IR(30) AND NOT IR(29) AND IR(28)) OR (IR(31) AND NOT IR(30) AND IR(29) AND NOT IR(28));
			MEM_READ <= IR(30);
			MEM_WRITE <= IR(29);
			WRITE_BACK <= IR(28);
			BRANCH <= IR(27) AND IR(26);
			JMP <= (IR(27) AND IR(26)) AND NOT(IR(25) OR IR(24) OR IR(23));
			HAS_NEXT_OPERAND <= IR(31);
			PUSH <= (NOT IR(27) AND IR(26) AND NOT IR(24) AND IR(25)) AND (NOT IR(23));
			POP <= (NOT IR(27) AND IR(26) AND NOT IR(24) AND IR(25)) AND (IR(23));

		END IF;
	END PROCESS;

END ARCHITECTURE;